`timescale 1ns / 1ps

module vga_controller(
    input wire clk_25mhz,       // 25 MHz clock
    input wire reset,           // Active high reset
    output wire hsync,          // Horizontal sync
    output wire vsync,          // Vertical sync
    output wire [9:0] h_count,  // Horizontal counter
    output wire [9:0] v_count,  // Vertical counter
    output wire display_enable  // High when in display area    
);

    // VGA 640x480 @ 60Hz timing parameters
    // Horizontal timing in pixels
    parameter H_DISPLAY = 640;      // Horizontal display width
    parameter H_FRONT   = 16;       // Front porch
    parameter H_SYNC    = 96;       // Sync pulse
    parameter H_BACK    = 48;       // Back porch
    parameter H_TOTAL   = H_DISPLAY + H_FRONT + H_SYNC + H_BACK; // Total cycle
    
    // Vertical timing in pixels
    parameter V_DISPLAY = 480;      // Vertical display height
    parameter V_FRONT   = 10;       // Front porch
    parameter V_SYNC    = 2;        // Sync pulse
    parameter V_BACK    = 33;       // Back porch
    parameter V_TOTAL   = V_DISPLAY + V_FRONT + V_SYNC + V_BACK; // Total cycle

endmodule
